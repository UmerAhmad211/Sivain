fun main() int {
	ret 0;	
}
